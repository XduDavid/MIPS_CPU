`include "defines.v"

module ex(
    input wire              rst,

    //����׶��͵�ִ�н׶ε���Ϣ
    input wire[`AluSelBus]  alusel_i,
    input wire[`AluOpBus]   aluop_i,
    input wire[`RegBus]     reg1_i,
    input wire[`RegBus]     reg2_i,
    input wire[`RegAddrBus] wd_i,
    input wire              wreg_i,

    //ִ�еĽ��
    output reg[`RegAddrBus] wd_o,       //ִ�н׶εĽ������Ҫд���Ŀ�ļĴ����ĵ�ַ
    output reg wreg_o,
    output reg[`RegBus] wdata_o,         //ִ�н׶�����Ҫд��Ŀ�ļĴ�����ֵ

    //����HI/LO����Ĵ�������ӵ��ź�
    input wire [31:0] hi_i,lo_i,    //HILOģ�������HI/LO�Ĵ�����ֵ
    //�ô�׶ε�����ǰ��
    input wire mem_whilo_i,         //���ڷô�׶ε�ָ���Ƿ�ҪдHI/LO�Ĵ���
    input wire [31:0] mem_hi_i,mem_lo_i, //���ڷô�׶ε�ָ��Ҫд��HI/LO�Ĵ�����ֵ
    //��д�׶ε�����ǰ��
    input wire wb_whilo_i,          //���ڻ�д�׶ε�ָ���Ƿ�Ҫд��HI/LO�Ĵ���
    input wire [31:0] wb_hi_i,wb_lo_i, //���ڻ�д�׶ε�ָ��Ҫд��HI/LO�Ĵ�����ֵ
    //HI/LO�����
    output reg whilo_o,
    output reg [31:0] hi_o,lo_o     //ִ�н׶ε�ָ��Ҫд��HI/LO�Ĵ�����ֵ
);

    //�����߼�����Ľ��
    reg [`RegBus] logicout;
    //������λ����Ľ��
    reg [`RegBus] shiftres;
    //�ƶ������Ľ��
    reg [`RegBus] moveres;

    //����HI/LO�Ĵ���������ֵ
    reg [`RegBus] HI,LO;

    //������������ı���
    reg[`RegBus] arithmeticres; //��������������
    wire ov_sum;				//����������
    wire reg1_eq_reg2;			//��һ���������Ƿ���ڵڶ���������
    wire reg1_lt_reg2;			//��һ���������Ƿ�С�ڵڶ���������
    wire[`RegBus] reg2_i_mux;	//��������ĵڶ�������reg2_i�Ĳ���
    wire[`RegBus] reg1_i_not;	//��������ĵ�һ��������reg1_iȡ�����ֵ
    wire[`RegBus] result_sum;	//����ӷ����
    wire[`RegBus] opdata1_mult;	//�˷������еı�����
    wire[`RegBus] opdata2_mult;	//�˷������еĳ���
    wire[`DoubleRegBus] hilo_temp;	//��ʱ����˷���������Ϊ64λ
    reg[`DoubleRegBus] mulres;		//����˷���������Ϊ64λ

//��������������ر�����ֵ
    //���Ϊ�������з��űȽ����㣬��reg2Ӧȡ������ʽ������ȡԭ��
    assign reg2_i_mux = ((aluop_i == `EXE_SUB_OP) || (aluop_i == `EXE_SUBU_OP) ||
                         (aluop_i == `EXE_SLT_OP)) ? (~reg2_i) + 1'b1 : reg2_i;
    //����Ǽӷ����㣬��reg2_i_mux=reg2_i������result_sum���Ǽӷ��Ľ��
    //����Ǽ������㣬��reg2_i_mux��reg2_i�Ĳ��룬����result_sum���Ǽ����Ľ��
    //������з��űȽ����㣬result_sum���Ǽ����Ľ�������ɸý����һ�����д�С���ж�
    assign result_sum = reg1_i + reg2_i_mux;
    //�Ӽ���ָ��ִ��ʱ�����жϽ���Ƿ���������������Ϊ���������������Ϊ����ʱ���������
    assign ov_sum = ((reg1_i[31] && reg2_i_mux[31] && (~result_sum[31]))) ||
                    (((~reg1_i[31] && ~reg2_i_mux[31]) && result_sum[31]));
    //�Ƚϲ�����1�Ƿ�С�ڲ�����2����з��űȽϺ��޷��űȽ����ַ�ʽ
    assign reg1_lt_reg2 = (aluop_i == `EXE_SLT_OP) ? ((reg1_i[31] && ~reg2_i[31]) ||
                          (~reg1_i[31] && ~reg2_i[31] && result_sum[31]) || 
                          (reg1_i[31] && reg2_i[31] && result_sum[31])): (reg1_i < reg2_i);
    //��reg_1��λȡ��������reg1_i_not
    assign reg1_i_not = ~reg1_i;
    //����1����Ϊ�з��ų˷��Ҹó���Ϊ��������ȡ�䲹�룬���򲻱�
    assign opdata1_mult = (((aluop_i == `EXE_MUL_OP) || (aluop_i == `EXE_MULT_OP))
                          && (reg1_i[31] == 1'b1)) ? (~reg1_i + 1'b1) : reg1_i;
    //����2����Ϊ�з��ų˷��Ҹó���Ϊ��������ȡ�䲹�룬���򲻱�
    assign opdata2_mult = (((aluop_i == `EXE_MUL_OP) || (aluop_i == `EXE_MULT_OP))
                          && (reg2_i[31] == 1'b1)) ? (~reg2_i + 1'b1) : reg2_i;
    //�õ���ʱ�ĳ˷���������浽hilo_temp��
    assign hilo_temp = opdata1_mult * opdata2_mult;
    //����ʱ�˷�������������������ս������mulres��
    always @(*) begin
        if(rst == `RstEnable) begin
            mulres = {`ZeroWord,`ZeroWord};
        end
        else if((aluop_i == `EXE_MUL_OP) || (aluop_i == `EXE_MULT_OP)) begin
            if(reg1_i[31] ^ reg2_i[31] == 1'b1) begin
                mulres = ~hilo_temp + 1'b1;
            end
            else begin
                mulres = hilo_temp;
            end
        end
        else begin
            mulres = hilo_temp;
        end
    end
/****************************************************
** �õ����µ�HI/LO�Ĵ�����ֵ���˴����������������   *****
****************************************************/
  always @(*) begin
    if(rst == `RstEnable) begin
      {HI,LO} <= {`ZeroWord,`ZeroWord};
    end
    else if(mem_whilo_i == `WriteEnable) begin
      {HI,LO} <= {mem_hi_i,mem_lo_i};
    end
    else if(wb_whilo_i == `WriteEnable) begin
      {HI,LO} <= {wb_hi_i,wb_lo_i};
    end
    else begin
      {HI,LO} <= {hi_i,lo_i};
    end
  end

/****************************************************
** MFHI��MFLO��MOVN��MOVZָ��(���дͨ�üĴ���������)  ***
****************************************************/
    always @(*) begin
      if(rst == `RstEnable) begin
          moveres = `ZeroWord;
      end
      else begin
          case(aluop_i)
              `EXE_MFHI_OP:   moveres = HI;
              `EXE_MFLO_OP:   moveres = LO;
              `EXE_MOVN_OP:   moveres = reg1_i;
              `EXE_MOVZ_OP:   moveres = reg1_i;
              default:        moveres = `ZeroWord;
          endcase
      end
    end


    //�����߼�����
    always @(*) begin
        if(rst == `RstEnable) begin
          logicout = `ZeroWord;
        end
        else begin
            case(aluop_i)
                `EXE_OR_OP:     logicout = reg1_i | reg2_i;
                `EXE_AND_OP:    logicout = reg1_i & reg2_i;
                `EXE_NOR_OP:    logicout = ~(reg1_i | reg2_i);
                `EXE_XOR_OP:    logicout = reg1_i ^ reg2_i;
                default:    logicout = `ZeroWord;
            endcase
        end  
    end

    //������λ����
    always @(*) begin
        if(rst == `RstEnable) begin
          shiftres = `ZeroWord;
        end
        else begin
          case(aluop_i)
            `EXE_SLL_OP:    shiftres = reg2_i << reg1_i[4:0];
            `EXE_SRL_OP:    shiftres = reg2_i >> reg1_i[4:0];
            `EXE_SRA_OP:begin
              shiftres = ({32{reg2_i[31]}}<<(6'd32-{1'b0,reg1_i[4:0]})) | (reg2_i >> reg1_i[4:0]);
            end
            default:        shiftres = `ZeroWord;
          endcase
        end
    end

    //������������
    always @(*) begin
        if(rst == `RstEnable) begin
            arithmeticres = `ZeroWord;
        end
        else begin
            case(aluop_i)
                `EXE_SLT_OP,`EXE_SLTU_OP:begin        //�Ƚ�����
                    arithmeticres = reg1_lt_reg2;
                end
                `EXE_ADD_OP,`EXE_ADDU_OP,`EXE_ADDI_OP,`EXE_ADDIU_OP:begin //�ӷ�����
                    arithmeticres = result_sum;
                end
                `EXE_SUB_OP,`EXE_SUBU_OP:begin        //��������
                    arithmeticres = result_sum;
                end
                `EXE_CLZ_OP:begin
                    arithmeticres = reg1_i[31] ? 0 : reg1_i[30] ? 1 : reg1_i[29] ? 2 :
													 reg1_i[28] ? 3 : reg1_i[27] ? 4 : reg1_i[26] ? 5 :
													 reg1_i[25] ? 6 : reg1_i[24] ? 7 : reg1_i[23] ? 8 : 
													 reg1_i[22] ? 9 : reg1_i[21] ? 10 : reg1_i[20] ? 11 :
													 reg1_i[19] ? 12 : reg1_i[18] ? 13 : reg1_i[17] ? 14 : 
													 reg1_i[16] ? 15 : reg1_i[15] ? 16 : reg1_i[14] ? 17 : 
													 reg1_i[13] ? 18 : reg1_i[12] ? 19 : reg1_i[11] ? 20 :
													 reg1_i[10] ? 21 : reg1_i[9] ? 22 : reg1_i[8] ? 23 : 
													 reg1_i[7] ? 24 : reg1_i[6] ? 25 : reg1_i[5] ? 26 : 
													 reg1_i[4] ? 27 : reg1_i[3] ? 28 : reg1_i[2] ? 29 : 
													 reg1_i[1] ? 30 : reg1_i[0] ? 31 : 32 ;
                end
                `EXE_CLO_OP:begin
                    arithmeticres = reg1_i_not[31] ? 0 : reg1_i_not[30] ? 1 : reg1_i_not[29] ? 2 :
													 reg1_i_not[28] ? 3 : reg1_i_not[27] ? 4 : reg1_i_not[26] ? 5 :
													 reg1_i_not[25] ? 6 : reg1_i_not[24] ? 7 : reg1_i_not[23] ? 8 : 
													 reg1_i_not[22] ? 9 : reg1_i_not[21] ? 10 : reg1_i_not[20] ? 11 :
													 reg1_i_not[19] ? 12 : reg1_i_not[18] ? 13 : reg1_i_not[17] ? 14 : 
													 reg1_i_not[16] ? 15 : reg1_i_not[15] ? 16 : reg1_i_not[14] ? 17 : 
													 reg1_i_not[13] ? 18 : reg1_i_not[12] ? 19 : reg1_i_not[11] ? 20 :
													 reg1_i_not[10] ? 21 : reg1_i_not[9] ? 22 : reg1_i_not[8] ? 23 : 
													 reg1_i_not[7] ? 24 : reg1_i_not[6] ? 25 : reg1_i_not[5] ? 26 : 
													 reg1_i_not[4] ? 27 : reg1_i_not[3] ? 28 : reg1_i_not[2] ? 29 : 
													 reg1_i_not[1] ? 30 : reg1_i_not[0] ? 31 : 32 ;
                end
                default:begin
                    arithmeticres = `ZeroWord;
                end
            endcase
        end
    end

    //�����MTHI��MTLOָ��������whilo_o,hi_o,lo_o��ֵ
    always @(*) begin
      if(rst == `RstEnable) begin
        whilo_o = `WriteDisable;
        hi_o = `ZeroWord;
        lo_o = `ZeroWord;
      end
      else if((aluop_i == `EXE_MULT_OP)||(aluop_i == `EXE_MULTU_OP)) begin
        whilo_o = `WriteEnable;
        hi_o = mulres[63:32];
        lo_o = mulres[31:0];
      end
      else if(aluop_i == `EXE_MTHI_OP) begin
        whilo_o = `WriteEnable;
        hi_o = reg1_i;
        lo_o = LO;        //дHI�Ĵ���������LO���ֲ���
      end
      else if(aluop_i == `EXE_MTLO_OP) begin
        whilo_o = `WriteEnable;
        hi_o = HI;        //дLO�Ĵ���������HI���ֲ���
        lo_o = reg1_i;        
      end
      else begin
        whilo_o = `WriteDisable;
        hi_o = `ZeroWord;
        lo_o = `ZeroWord;
      end
    end

    //����aluselָʾ���������ͣ�ѡ��һ����������Ϊ���ս��
    //��ʱֻ���߼�������
    always @(*) begin
        wd_o = wd_i;
          if(((aluop_i == `EXE_ADD_OP) || (aluop_i == `EXE_ADDI_OP) || 
            (aluop_i == `EXE_SUB_OP)) && (ov_sum == 1'b1))begin
              wreg_o = `WriteDisable;
          end
          else begin
              wreg_o = wreg_i;
          end
        case(alusel_i)
            `EXE_RES_LOGIC:     wdata_o = logicout;
            `EXE_RES_SHIFT:     wdata_o = shiftres;
            `EXE_RES_MOVE:      wdata_o = moveres;
            `EXE_RES_ARITHMETIC:wdata_o = arithmeticres;
            `EXE_RES_MUL:       wdata_o = mulres;
            default:            wdata_o = `ZeroWord;
        endcase
    end

endmodule